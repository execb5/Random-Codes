
library ieee ;
	use ieee.std_logic_1164.all ;
	use ieee.numeric_std.all ;

entity SodaMachine is
	port(
			M025, M050, M100, DEV, SUCO, AGUA, reset, ck : in std_logic;
			D025, D050, D100, L_SUCO, L_AGUA, insuficienteOut : out std_logic;
			centena, dezena, unidade : out std_logic_vector(3 downto 0)
		);
end entity ; -- SodaMachine

architecture Behavioral of SodaMachine is
	type myDearStates is (R0_00, R0_25, R0_50, R0_75, R1_00, R1_25, R1_50, R1_75);
	signal currentState : myDearStates;
	signal insuficiente : std_logic;
begin

	insuficienteOut <= insuficiente;

	process(ck)
	begin
		if (ck'event and ck = '1') then
			centena <= "0000";
			dezena <= "0000";
			unidade <= "0000";
			insuficiente <= '0';
			D025 <= '0';
			D050 <= '0';
			D100 <= '0';
			L_AGUA <= '0';
			L_SUCO <= '0';
			if (reset = '1') then
				currentState <= R0_00;
				centena <= "0000";
				dezena <= "0000";
				unidade <= "0000";
				insuficiente <= '0';
				D025 <= '0';
				D050 <= '0';
				D100 <= '0';
				L_AGUA <= '0';
				L_SUCO <= '0';
			else
				case(currentState) is
					when R0_00 =>
						if (M025 = '1') then
							currentState <= R0_25;
							centena <= "0000";
							dezena <= "0010";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M050 = '1') then
							currentState <= R0_50;
							centena <= "0000";
							dezena <= "0101";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M100 = '1') then
							currentState <= R1_00;
							centena <= "0001";
							dezena <= "0000";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (DEV = '1') then
							currentState <= R0_00;
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (SUCO = '1') then
							insuficiente <= '1';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (AGUA = '1') then
							insuficiente <= '1';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						end if ;
					when R0_25 =>
						if (M025 = '1') then
							currentState <= R0_50;
							centena <= "0000";
							dezena <= "0101";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M050 = '1') then
							currentState <= R0_75;
							centena <= "0000";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M100 = '1') then
							currentState <= R1_25;
							centena <= "0001";
							dezena <= "0010";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (DEV = '1') then
							currentState <= R0_00;
							centena <= "0000";
							dezena <= "0000";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (SUCO = '1') then
							insuficiente <= '1';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (AGUA = '1') then
							insuficiente <= '1';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						end if ;
					when R0_50 =>
						if (M025 = '1') then
							currentState <= R0_75;
							centena <= "0000";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M050 = '1') then
							currentState <= R1_00;
							centena <= "0001";
							dezena <= "0000";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M100 = '1') then
							currentState <= R1_50;
							centena <= "0001";
							dezena <= "0101";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (DEV = '1') then
							currentState <= R0_00;
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '1';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (SUCO = '1') then
							insuficiente <= '1';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (AGUA = '1') then
							insuficiente <= '1';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						end if ;
					when R0_75 =>
						if (M025 = '1') then
							currentState <= R1_00;
							centena <= "0001";
							dezena <= "0000";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M050 = '1') then
							currentState <= R1_25;
							centena <= "0001";
							dezena <= "0010";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M100 = '1') then
							currentState <= R1_75;
							centena <= "0001";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (DEV = '1') then
							currentState <= R0_00;
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '1';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (SUCO = '1') then
							insuficiente <= '1';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (AGUA = '1') then
							insuficiente <= '1';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						end if ;
					when R1_00 =>
						if (M025 = '1') then
							currentState <= R1_25;
							centena <= "0001";
							dezena <= "0010";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M050 = '1') then
							currentState <= R1_50;
							centena <= "0001";
							dezena <= "0101";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M100 = '1') then
							currentState <= R1_75;
							centena <= "0001";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (DEV = '1') then
							currentState <= R0_00;
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '1';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (SUCO = '1') then
							insuficiente <= '1';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (AGUA = '1') then
							currentState <= R0_00;
							centena <= "0000";
							dezena <= "0000";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '1';
							L_SUCO <= '0';
						end if;
					when R1_25 =>
						if (M025 = '1') then
							currentState <= R1_50;
							centena <= "0001";
							dezena <= "0101";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M050 = '1') then
							currentState <= R1_75;
							centena <= "0001";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M100 = '1') then
							currentState <= R1_75;
							centena <= "0001";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '1';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (DEV = '1') then
							currentState <= R0_00;
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '0';
							D100 <= '1';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (SUCO = '1') then
							insuficiente <= '1';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (AGUA = '1') then
							currentState <= R0_00;
							centena <= "0000";
							dezena <= "0000";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '1';
							L_SUCO <= '0';
						end if;
					when R1_50 =>
						if (M025 = '1') then
							currentState <= R1_75;
							centena <= "0001";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M050 = '1') then
							currentState <= R1_75;
							centena <= "0001";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M100 = '1') then
							currentState <= R1_75;
							centena <= "0001";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '1';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (DEV = '1') then
							currentState <= R0_00;
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '1';
							D100 <= '1';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (SUCO = '1') then
							currentState <= R0_00;
							centena <= "0000";
							dezena <= "0000";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '1';
						elsif (AGUA = '1') then
							currentState <= R0_00;
							centena <= "0000";
							dezena <= "0000";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '1';
							D100 <= '0';
							L_AGUA <= '1';
							L_SUCO <= '0';
						end if;
					when R1_75 =>
						if (M025 = '1') then
							currentState <= R1_75;
							centena <= "0001";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M050 = '1') then
							currentState <= R1_75;
							centena <= "0001";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '1';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (M100 = '1') then
							currentState <= R1_75;
							centena <= "0001";
							dezena <= "0111";
							unidade <= "0101";
							insuficiente <= '0';
							D025 <= '0';
							D050 <= '0';
							D100 <= '1';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (DEV = '1') then
							currentState <= R0_00;
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '1';
							D100 <= '1';
							L_AGUA <= '0';
							L_SUCO <= '0';
						elsif (SUCO = '1') then
							currentState <= R0_00;
							centena <= "0000";
							dezena <= "0000";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '0';
							D100 <= '0';
							L_AGUA <= '0';
							L_SUCO <= '1';
						elsif (AGUA = '1') then
							currentState <= R0_00;
							centena <= "0000";
							dezena <= "0000";
							unidade <= "0000";
							insuficiente <= '0';
							D025 <= '1';
							D050 <= '1';
							D100 <= '0';
							L_AGUA <= '1';
							L_SUCO <= '0';
						end if ;
				end case ;
			end if ;
		end if ;
	end process ;
end architecture ; -- Behavioral